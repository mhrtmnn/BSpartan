package AxiBridge;

import ClientServer::*;
import GlobalTypes::*;
import GetPut::*;
import FIFO::*;


/******************************************************
* GLOBAL TYPES/FUNCTIONS/DATA
******************************************************/
typedef enum { NVALID, VALID } AxiValid deriving (Bits);

typedef enum {
	OKAY,	// Normal access okay
	EXOKAY,	// Exclusive access okay
	SLVERR,	// Access has reached the slave okay, but slave wishes to indicate error condition
	DECERR	// Typically generated by an interconnect to indicate that there is no slave at the address
} AxiRespCode deriving (Bits, Eq, FShow);

typedef struct {
	Bit#(a_len) 			addr;
	Bit#(TDiv#(d_len, 8)) 	strobe;
	Bit#(d_len) 			data;
} AXI_TX_tfer#(numeric type d_len, numeric type a_len) deriving (Bits);

typedef struct {
	Bit#(a_len) 			addr;
} AXI_RX_tfer#(numeric type a_len) deriving (Bits);

// helper function TX
function Action axilite_send(AxiBridge#(d, a) axi, Bit#(a) addr, Bit#(n) data) provisos(Add#(n, _unused, d));
action
	let t = AXI_TX_tfer {
		addr 	: addr,
		data 	: extend(data),
		strobe 	: fromInteger(get_strobe(data))
	};
	axi.tx.put(t);
endaction
endfunction

// helper function RX 1
function Action axilite_recv_start(AxiBridge#(d, a) axi, Bit#(a) addr);
action
	let t = AXI_RX_tfer {
		addr:addr
	};
	axi.rx.request.put(t);
endaction
endfunction

// helper function RX 2
function ActionValue#(Bit#(d)) axilite_recv_get(AxiBridge#(d, a) axi);
actionvalue
	let val <- axi.rx.response.get();
	return val;
endactionvalue
endfunction


/******************************************************
* FUNCTIONS
******************************************************/
function Integer get_strobe(Bit#(sz) b);
	return valueOf(TDiv#(sz, 8));
endfunction


/******************************************************
* GENERIC AXI IFACE
******************************************************/
interface AxiLiteIface#(numeric type d_len, numeric type a_len);
	method Action putCLK(bit clk);

	// AW Channel
	method Action putAW(Bit#(a_len) awaddr, bit awvalid);
	method bit getAWready();

	// W Channel
	method Action putW(Bit#(d_len) wdata, bit wvalid, Bit#(TDiv#(d_len, 8)) wstrb);
	method bit getWready();

	// B Channel
	method Action putB(bit bready);
	method bit getBvalid();
	method Bit#(2) getBresp();

	// AR Channel
	method Action putAR(Bit#(a_len) araddr, bit arvalid);
	method bit getARready();

	// R Channel
	method Action putR(bit rready);
	method bit getRvalid();
	method Bit#(d_len) getRdata();
	method Bit#(2) getRresp();
endinterface


/******************************************************
* BSV AXI INTERFACE
******************************************************/
interface AxiBridge#(numeric type d_len, numeric type a_len);
	interface Server#(AXI_RX_tfer#(a_len), Bit#(d_len)) 	rx;
	interface Put#(AXI_TX_tfer#(d_len, a_len)) 				tx;
endinterface

module mkAxiBridge#(AxiLiteIface#(d_len, a_len) coreAXI) (AxiBridge#(d_len, a_len))
	provisos (Div#(d_len, 8, stb_len));

	/* RX iface */
	FIFO#(AXI_RX_tfer#(a_len)) 			rx_fifo_in		<- mkFIFO();
	FIFO#(Bit#(d_len)) 					rx_fifo_out		<- mkFIFO();

	Reg#(Bool) 							pending_r_addr 	<- mkReg(True);

	/* TX iface */
	FIFO#(AXI_TX_tfer#(d_len, a_len)) 	tx_fifo_in		<- mkFIFO();

	Reg#(Bool) 							pending_w_addr 	<- mkReg(True);
	Reg#(Bool) 							pending_w_data 	<- mkReg(True);

	/* module state */
	Reg#(bit) clk 					<- mkReg(0);
	Reg#(Int#(4)) axi_w_state 		<- mkReg(0);
	Reg#(Int#(4)) axi_aw_state 		<- mkReg(0);
	Reg#(Int#(4)) axi_r_state 		<- mkReg(0);
	Reg#(Int#(4)) axi_ar_state 		<- mkReg(0);

	/* buffer for axi signals */
	Reg#(Bit#(  a_len)) buf_awaddr 	<- mkReg(0);
	Reg#(Bit#(      1)) buf_awvalid	<- mkReg(0);
	Reg#(Bit#(  d_len)) buf_wdata 	<- mkReg(0);
	Reg#(Bit#(      1)) buf_wvalid 	<- mkReg(0);
	Reg#(Bit#(stb_len)) buf_wstrb 	<- mkReg(0);
	Reg#(Bit#(      1)) buf_bready 	<- mkReg(0);
	Reg#(Bit#(  a_len)) buf_araddr	<- mkReg(0);
	Reg#(Bit#(      1)) buf_arvalid	<- mkReg(0);
	Reg#(Bit#(      1)) buf_rready 	<- mkReg(0);


	/******************************************************
	* RULES
	******************************************************/


	/******************** IFACE RULES ********************/

	rule axi_tx_iface(!pending_w_addr && !pending_w_data);
		$display("[AXIlite] [%d] Deq from tx_fifo_in", $time);

		// discard head, which was successfully transferred
		tx_fifo_in.deq();

		pending_w_addr <= True;
		pending_w_data <= True;
	endrule

	rule axi_rx_iface(!pending_r_addr);
		$display("[AXIlite] [%d] Deq from rx_fifo_in", $time);

		// discard head, which was successfully transferred
		rx_fifo_in.deq();

		pending_r_addr <= True;
	endrule


	/********************** AXI READ *********************/

	// R Channel
	rule axi_R(clk == 1 && axi_r_state == 0);
		let r_resp 	= coreAXI.getRresp();
		let r_valid = coreAXI.getRvalid();

		// rule only fires if FIFO is not full, ie wen can receive data
		buf_rready 	<= 1;

		if (r_valid == pack(VALID) && r_resp == pack(OKAY)) begin

			// read data
			let r_data 	= coreAXI.getRdata();
			rx_fifo_out.enq(r_data);

			axi_r_state <= 1;
		end
	endrule

	rule axi_R_idle(clk == 1 && axi_r_state == 1);
		buf_rready 	<= 0;
		axi_r_state <= 0;
	endrule


	// AR Channel
	rule axi_AR(clk == 1 && pending_r_addr && axi_ar_state == 0);

		// change signal levels once clock goes low
		buf_araddr 		<= rx_fifo_in.first.addr;
		buf_arvalid 	<= pack(VALID);

		axi_ar_state 	<= 1;
	endrule

	rule axi_AR_ctrl(clk == 1 && pending_r_addr && axi_ar_state == 1);

		// read signal levels while clock is high
		if (coreAXI.getARready() == 1) begin
			axi_ar_state <= 2;
		end
	endrule

	rule axi_AR_ctrl1(clk == 1 && pending_r_addr && axi_ar_state == 2);

		// change signal levels once clock goes low
		buf_araddr  	<= 0;
		buf_arvalid 	<= pack(NVALID);

		pending_r_addr 	<= False;
		axi_ar_state 	<= 0;
	endrule


	/********************** AXI WRITE ********************/

	// AW Channel
	rule axi_AW(clk == 1 && pending_w_addr && axi_aw_state == 0);

		// change signal levels once clock goes low
		buf_awaddr 		<= tx_fifo_in.first.addr;
		buf_awvalid 	<= pack(VALID);

		axi_aw_state 	<= 1;
	endrule

	rule axi_AW_ctrl(clk == 1 && pending_w_addr && axi_aw_state == 1);

		// read signal levels while clock is high
		if (coreAXI.getAWready() == 1) begin
			axi_aw_state <= 2;
		end
	endrule

	rule axi_AW_ctrl1(clk == 1 && pending_w_addr && axi_aw_state == 2);

		// change signal levels once clock goes low
		buf_awaddr 		<= 0;
		buf_awvalid 	<= pack(NVALID);

		// synchronize Channel AW and W in tule axi_B
	endrule

	// W Channel
	rule axi_W(clk == 1 && pending_w_data && axi_w_state == 0);

		// change signal levels once clock goes low
		buf_wdata 	<= tx_fifo_in.first.data;
		buf_wstrb 	<= tx_fifo_in.first.strobe;
		buf_wvalid 	<= pack(VALID);

		axi_w_state <= 1;
	endrule

	rule axi_W_ctrl(clk == 1 && pending_w_data && axi_w_state == 1);

		// read signal levels while clock is high
		if (coreAXI.getWready() == 1) begin
			axi_w_state <= 2;
		end
	endrule

	rule axi_W_ctrl1(clk == 1 && pending_w_data && axi_w_state == 2);

		// change signal levels once clock goes low
		buf_wdata 	<= 0;
		buf_wstrb 	<= 0;
		buf_wvalid 	<= pack(NVALID);

		// synchronize Channel AW and W in tule axi_B
	endrule

	// B Channel
	rule axi_B(clk == 1 && axi_w_state == 2 && axi_aw_state == 2 && pending_w_data && pending_w_addr);

		// always ready to receive
		buf_bready 	<= 1;

		let b_valid = coreAXI.getBvalid();
		let b_resp  = coreAXI.getBresp();

		if (b_valid == pack(VALID)) begin
			if (b_resp == pack(OKAY)) begin
				pending_w_addr <= False;
				pending_w_data <= False;
			end else begin
				$display("[AXIlite] AXI Write Error: %d (retrying)", b_resp);
			end

			axi_w_state 	<= 0;
			axi_aw_state 	<= 0;
		end
	endrule


	/*********************** SYSTEM **********************/

	rule axi_clk;
		clk <= ~clk;
		coreAXI.putCLK(clk);
	endrule

	/* drive signals in every cycle */
	(*fire_when_enabled*)
	rule signal_driver;
		coreAXI.putAW(buf_awaddr, buf_awvalid);
		coreAXI.putW(buf_wdata, buf_wvalid, buf_wstrb);
		coreAXI.putB(buf_bready);
		coreAXI.putAR(buf_araddr, buf_arvalid);
		coreAXI.putR(buf_rready);
	endrule


	/******************************************************
	* INTERFACE
	******************************************************/
	interface Server rx;
		interface Put request 	= toPut(rx_fifo_in);
		interface Get response 	= toGet(rx_fifo_out);
	endinterface

	interface tx = toPut(tx_fifo_in);

endmodule

endpackage
