package GlobalTypes;


/******************************************************
* GLOBAL TYPES/FUNCTIONS/DATA
******************************************************/
typedef Bit#(8) Byte;

endpackage
